module fulladder(
input A,
input B,
input C_IN,
output C_OUT,
output S);
c_addsub_0 fa(.A(A),.B(B),.C_IN(C_IN),.C_OUT(C_OUT),.S(S));
endmodule
